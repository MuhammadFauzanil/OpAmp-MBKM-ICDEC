magic
tech sky130A
magscale 1 2
timestamp 1729217204
<< nwell >>
rect -176 -690 822 2170
<< nsubdiff >>
rect -140 2100 -80 2134
rect 726 2100 786 2134
rect -140 2074 -106 2100
rect 752 2074 786 2100
rect -140 -620 -106 -594
rect 752 -620 786 -594
rect -140 -654 -80 -620
rect 726 -654 786 -620
<< nsubdiffcont >>
rect -80 2100 726 2134
rect -140 -594 -106 2074
rect 752 -594 786 2074
rect -80 -654 726 -620
<< poly >>
rect -56 2062 36 2078
rect -56 2028 -40 2062
rect -6 2028 36 2062
rect -56 2012 36 2028
rect 6 1981 36 2012
rect 610 2062 702 2078
rect 610 2028 652 2062
rect 686 2028 702 2062
rect 610 2012 702 2028
rect 610 2004 640 2012
rect -56 1368 36 1384
rect 94 1383 294 1485
rect -56 1334 -40 1368
rect -6 1334 36 1368
rect -56 1318 36 1334
rect 6 1287 36 1318
rect 610 1368 702 1384
rect 610 1334 652 1368
rect 686 1334 702 1368
rect 610 1318 702 1334
rect 610 1287 640 1318
rect 94 690 552 790
rect 6 162 36 193
rect -56 146 36 162
rect -56 112 -40 146
rect -6 112 36 146
rect -56 96 36 112
rect 610 162 640 193
rect 610 146 702 162
rect 610 112 652 146
rect 686 112 702 146
rect 610 96 702 112
rect 352 -4 552 96
rect 6 -532 36 -501
rect -56 -548 36 -532
rect -56 -582 -40 -548
rect -6 -582 36 -548
rect -56 -598 36 -582
rect 610 -532 640 -501
rect 610 -548 702 -532
rect 610 -582 652 -548
rect 686 -582 702 -548
rect 610 -598 702 -582
<< polycont >>
rect -40 2028 -6 2062
rect 652 2028 686 2062
rect -40 1334 -6 1368
rect 652 1334 686 1368
rect -40 112 -6 146
rect 652 112 686 146
rect -40 -582 -6 -548
rect 652 -582 686 -548
<< locali >>
rect -140 2100 -80 2134
rect 726 2100 786 2134
rect -140 2074 -106 2100
rect 752 2074 786 2100
rect -56 2028 -40 2062
rect -6 2028 10 2062
rect 636 2028 652 2062
rect 686 2028 702 2062
rect -40 1981 -6 2028
rect 652 1975 686 2028
rect -56 1334 -40 1368
rect -6 1334 10 1368
rect 636 1334 652 1368
rect 686 1334 702 1368
rect -40 1287 -6 1334
rect 652 1287 686 1334
rect -40 146 -6 193
rect 652 146 686 193
rect -56 112 -40 146
rect -6 112 10 146
rect 636 112 652 146
rect 686 112 702 146
rect -40 -548 -6 -501
rect 652 -548 686 -501
rect -56 -582 -40 -548
rect -6 -582 10 -548
rect 636 -582 652 -548
rect 686 -582 702 -548
rect -140 -620 -106 -594
rect 752 -620 786 -594
rect -140 -654 -80 -620
rect 726 -654 786 -620
<< viali >>
rect 652 2100 686 2134
rect -40 2028 -6 2062
rect 652 2028 686 2062
rect -40 1334 -6 1368
rect 652 1334 686 1368
rect -40 112 -6 146
rect 652 112 686 146
rect -40 -582 -6 -548
rect 652 -582 686 -548
rect -40 -654 -6 -620
<< metal1 >>
rect 640 2134 698 2140
rect 640 2100 652 2134
rect 686 2100 698 2134
rect -52 2062 6 2068
rect -52 2028 -40 2062
rect -6 2028 6 2062
rect -52 2022 6 2028
rect 640 2062 698 2100
rect 640 2028 652 2062
rect 686 2028 698 2062
rect 640 2022 698 2028
rect -47 1981 0 2022
rect 646 1981 693 2022
rect -47 1969 88 1981
rect -59 1593 -49 1969
rect 3 1593 88 1969
rect -46 1581 88 1593
rect 300 1540 346 1981
rect 558 1968 693 1981
rect 558 1581 692 1968
rect 558 1540 604 1581
rect 300 1494 604 1540
rect -52 1368 6 1374
rect -52 1334 -40 1368
rect -6 1334 6 1368
rect -52 1328 6 1334
rect -47 1287 0 1328
rect -40 1276 94 1287
rect -40 1275 101 1276
rect -40 899 39 1275
rect 91 899 101 1275
rect -40 887 94 899
rect 42 634 134 680
rect 42 593 88 634
rect -46 193 88 593
rect -47 152 0 193
rect -52 146 6 152
rect -52 112 -40 146
rect -6 112 6 146
rect -52 106 6 112
rect 300 -13 346 1494
rect 640 1368 698 1374
rect 640 1334 652 1368
rect 686 1334 698 1368
rect 640 1328 698 1334
rect 646 1287 693 1328
rect 558 911 692 1287
rect 557 887 692 911
rect 557 846 603 887
rect 515 800 603 846
rect 558 582 692 593
rect 545 205 555 582
rect 607 205 692 582
rect 558 193 692 205
rect 646 152 693 193
rect 640 146 698 152
rect 640 112 652 146
rect 686 112 698 146
rect 640 106 698 112
rect 42 -59 346 -13
rect 42 -101 88 -59
rect -47 -109 88 -101
rect -47 -110 87 -109
rect -47 -501 88 -110
rect 300 -501 346 -59
rect 552 -113 688 -101
rect 552 -489 643 -113
rect 695 -489 705 -113
rect 552 -501 693 -489
rect -47 -542 0 -501
rect 646 -542 693 -501
rect -52 -548 6 -542
rect -52 -582 -40 -548
rect -6 -582 6 -548
rect -52 -620 6 -582
rect 640 -548 698 -542
rect 640 -582 652 -548
rect 686 -582 698 -548
rect 640 -588 698 -582
rect -52 -654 -40 -620
rect -6 -654 6 -620
rect -52 -660 6 -654
<< via1 >>
rect -49 1593 3 1969
rect 39 899 91 1275
rect 555 205 607 582
rect 643 -489 695 -113
<< metal2 >>
rect -49 1969 3 1979
rect -49 1472 3 1593
rect -58 1462 3 1472
rect 639 1462 699 1472
rect 2 1402 3 1462
rect 630 1402 639 1462
rect 699 1402 708 1462
rect -58 1392 3 1402
rect 639 1392 699 1402
rect -49 83 3 1392
rect 39 1275 91 1285
rect 91 899 92 912
rect 39 889 92 899
rect 40 767 92 889
rect 40 715 607 767
rect 555 582 607 715
rect 555 195 607 205
rect 643 83 695 1392
rect -53 73 7 83
rect 641 73 701 83
rect -62 13 -53 73
rect 7 13 16 73
rect -53 3 7 13
rect 641 3 701 13
rect 643 -113 695 3
rect 643 -499 695 -489
<< via2 >>
rect -58 1402 2 1462
rect 639 1402 699 1462
rect -53 13 7 73
rect 641 13 701 73
<< metal3 >>
rect -68 1462 12 1467
rect 629 1462 709 1467
rect -68 1402 -58 1462
rect 2 1402 639 1462
rect 699 1402 709 1462
rect -68 1397 12 1402
rect 629 1397 709 1402
rect -63 73 17 78
rect 631 73 711 78
rect -63 13 -53 73
rect 7 13 641 73
rect 701 13 711 73
rect -63 8 17 13
rect 631 8 711 13
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_0
timestamp 1729134163
transform 1 0 21 0 1 1087
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_1
timestamp 1729134163
transform 1 0 21 0 1 -301
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_2
timestamp 1729134163
transform 1 0 625 0 1 -301
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_3
timestamp 1729134163
transform 1 0 625 0 1 393
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_4
timestamp 1729134163
transform 1 0 21 0 1 393
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_5
timestamp 1729134163
transform 1 0 625 0 1 1087
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_6
timestamp 1729134163
transform 1 0 21 0 1 1781
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_2ZH9AN  sky130_fd_pr__pfet_01v8_2ZH9AN_7
timestamp 1729134163
transform 1 0 625 0 1 1781
box -109 -262 109 262
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_0
timestamp 1729141650
transform 1 0 323 0 1 1781
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_1
timestamp 1729141650
transform 1 0 323 0 1 1087
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_2
timestamp 1729141650
transform 1 0 323 0 1 393
box -323 -300 323 300
use sky130_fd_pr__pfet_01v8_SDE6B7  sky130_fd_pr__pfet_01v8_SDE6B7_3
timestamp 1729141650
transform 1 0 323 0 1 -301
box -323 -300 323 300
<< labels >>
flabel metal1 s 666 2076 666 2076 0 FreeSans 1600 0 0 0 VDD
port 0 nsew
flabel metal2 s 56 812 56 812 0 FreeSans 1600 0 0 0 D1
port 1 nsew
flabel metal1 s 580 842 580 842 0 FreeSans 1600 0 0 0 D2
port 2 nsew
flabel metal3 s 534 1434 534 1434 0 FreeSans 1600 0 0 0 D5
port 3 nsew
<< end >>
