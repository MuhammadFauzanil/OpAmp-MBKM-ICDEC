magic
tech sky130A
magscale 1 2
timestamp 1729356413
<< nwell >>
rect 845 -2214 1250 -1412
<< viali >>
rect 2252 -825 2286 -791
rect 1758 -977 1823 -941
rect 1170 -1278 1514 -1044
rect 1590 -1278 1934 -1044
rect 2004 -1279 2348 -1045
rect 3244 -1280 3588 -1046
<< metal1 >>
rect 2236 -791 2379 -778
rect 1746 -941 1835 -935
rect 1746 -977 1758 -941
rect 1823 -977 1835 -941
rect 1746 -1038 1835 -977
rect 1158 -1044 1526 -1038
rect 1158 -1162 1170 -1044
rect 988 -1207 1170 -1162
rect 114 -2157 159 -2099
rect 988 -2157 1033 -1207
rect 1158 -1278 1170 -1207
rect 1514 -1278 1526 -1044
rect 1158 -1284 1526 -1278
rect 1578 -1044 1946 -1038
rect 2158 -1039 2200 -793
rect 2236 -825 2252 -791
rect 2286 -825 2379 -791
rect 2236 -836 2379 -825
rect 2321 -844 2379 -836
rect 3044 -844 3102 -809
rect 2321 -902 3102 -844
rect 1578 -1278 1590 -1044
rect 1934 -1278 1946 -1044
rect 1578 -1284 1946 -1278
rect 1992 -1045 2360 -1039
rect 1992 -1279 2004 -1045
rect 2348 -1279 2360 -1045
rect 3232 -1046 3600 -1040
rect 1992 -1285 2360 -1279
rect 2434 -1280 2444 -1046
rect 2788 -1280 2798 -1046
rect 2840 -1280 2850 -1046
rect 3194 -1280 3204 -1046
rect 3232 -1280 3244 -1046
rect 3588 -1280 3600 -1046
rect 2158 -1364 2200 -1285
rect 3232 -1286 3600 -1280
rect 3394 -1354 3436 -1286
rect 1227 -1406 2200 -1364
rect 1227 -1740 1269 -1406
rect 2649 -1425 2659 -1373
rect 2779 -1425 2799 -1373
rect 2766 -1694 2799 -1425
rect 2842 -1396 3436 -1354
rect 2842 -1723 2884 -1396
rect 114 -2202 1033 -2157
<< via1 >>
rect 2444 -1280 2788 -1046
rect 2850 -1280 3194 -1046
rect 2659 -1425 2779 -1373
<< metal2 >>
rect 1660 -978 1712 -788
rect 2936 -821 2982 -637
rect 1084 -1030 1712 -978
rect 2601 -867 2982 -821
rect 1084 -1294 1136 -1030
rect 2601 -1036 2647 -867
rect 2444 -1046 2788 -1036
rect 2444 -1290 2788 -1280
rect 2850 -1046 3194 -1036
rect 2850 -1290 3194 -1280
rect 1084 -1346 1791 -1294
rect 2966 -1318 3019 -1290
rect 1739 -1582 1791 -1346
rect 2659 -1371 3019 -1318
rect 2659 -1373 2779 -1371
rect 2659 -1435 2779 -1425
<< metal3 >>
rect 789 -1510 1043 -1449
rect 982 -1782 1043 -1510
rect 982 -1843 1633 -1782
use nmos_dif  nmos_dif_0
timestamp 1729345511
transform 0 1 1266 -1 0 473
box -176 -198 1448 1019
use nmosrs  nmosrs_0
timestamp 1729225292
transform 1 0 2673 0 1 -1
box -292 -819 978 647
use pmos_dif  pmos_dif_0
timestamp 1729246480
transform 0 1 2419 -1 0 -1590
box -176 -1316 622 1231
use pmoscs  pmoscs_0
timestamp 1729217204
transform 1 0 160 0 1 -1522
box -176 -690 822 2170
<< labels >>
flabel via1 3016 -1171 3016 -1171 0 FreeSans 480 0 0 0 VIN
port 4 nsew
flabel viali 3416 -1173 3416 -1173 0 FreeSans 480 0 0 0 VIP
port 5 nsew
flabel via1 2624 -1172 2624 -1172 0 FreeSans 480 0 0 0 RS
port 3 nsew
flabel viali 2189 -1172 2189 -1172 0 FreeSans 480 0 0 0 OUT
port 2 nsew
flabel viali 1757 -1173 1757 -1173 0 FreeSans 480 0 0 0 GND
port 1 nsew
flabel viali 1339 -1173 1339 -1173 0 FreeSans 480 0 0 0 VDD
port 0 nsew
<< end >>
