magic
tech sky130A
magscale 1 2
timestamp 1729345511
<< psubdiff >>
rect -176 985 -90 1019
rect 1385 985 1448 1019
rect -176 959 -142 985
rect 1414 959 1448 985
rect -176 -146 -142 -120
rect 1414 -146 1448 -120
rect -176 -180 -87 -146
rect 1388 -180 1448 -146
<< psubdiffcont >>
rect -90 985 1385 1019
rect -176 -120 -142 959
rect 1414 -120 1448 959
rect -87 -180 1388 -146
<< poly >>
rect -30 524 0 532
rect -92 508 0 524
rect -92 474 -76 508
rect -42 474 0 508
rect -92 458 0 474
rect 1272 523 1302 558
rect 1272 507 1364 523
rect 1272 473 1314 507
rect 1348 473 1364 507
rect 1272 457 1364 473
rect -92 372 0 388
rect -92 338 -76 372
rect -42 338 0 372
rect -92 322 0 338
rect -30 314 0 322
rect 1272 372 1364 388
rect 1272 338 1314 372
rect 1348 338 1364 372
rect 1272 322 1364 338
rect 1272 314 1302 322
<< polycont >>
rect -76 474 -42 508
rect 1314 473 1348 507
rect -76 338 -42 372
rect 1314 338 1348 372
<< locali >>
rect -176 985 -90 1019
rect 1385 985 1448 1019
rect -176 959 -142 985
rect 1414 959 1448 985
rect -76 508 -42 562
rect -92 474 -76 508
rect -42 474 -26 508
rect 1314 507 1348 563
rect 1298 473 1314 507
rect 1348 473 1364 507
rect -92 338 -76 372
rect -42 338 -26 372
rect 1298 338 1314 372
rect 1348 338 1364 372
rect -76 282 -42 338
rect 1313 282 1348 338
rect -176 -146 -142 -120
rect 1414 -146 1448 -120
rect -176 -180 -87 -146
rect 1388 -180 1448 -146
<< viali >>
rect -76 474 -42 508
rect 1314 473 1348 507
rect -76 338 -42 372
rect 1314 338 1348 372
rect 933 -146 998 -144
rect 277 -180 329 -146
rect 933 -180 998 -146
rect 933 -181 998 -180
<< metal1 >>
rect 604 936 610 941
rect -36 894 610 936
rect -36 758 6 894
rect 604 889 610 894
rect 662 936 668 941
rect 662 894 1308 936
rect 662 889 668 894
rect 1266 758 1308 894
rect -82 558 52 758
rect 224 558 384 758
rect 556 558 716 758
rect 888 558 1048 758
rect 1220 558 1354 758
rect -82 514 -36 558
rect -88 508 -30 514
rect -88 474 -76 508
rect -42 474 -30 508
rect 64 477 74 529
rect 202 477 212 529
rect -88 468 -30 474
rect -88 372 -30 378
rect -88 338 -76 372
rect -42 338 -30 372
rect -88 332 -30 338
rect -82 288 -36 332
rect 64 317 74 369
rect 202 317 212 369
rect 275 288 331 558
rect 610 529 662 558
rect 600 520 610 529
rect 540 486 610 520
rect 600 477 610 486
rect 662 520 672 529
rect 662 486 735 520
rect 662 477 672 486
rect 396 317 406 369
rect 534 317 544 369
rect 728 317 738 369
rect 866 317 876 369
rect 940 288 996 558
rect 1060 477 1070 529
rect 1198 477 1208 529
rect 1308 513 1354 558
rect 1302 507 1360 513
rect 1302 473 1314 507
rect 1348 473 1360 507
rect 1302 467 1360 473
rect 1302 372 1360 378
rect 1060 317 1070 369
rect 1198 317 1208 369
rect 1302 338 1314 372
rect 1348 338 1360 372
rect 1302 332 1360 338
rect 1307 289 1354 332
rect -82 276 52 288
rect -82 100 -41 276
rect 11 100 52 276
rect -82 88 52 100
rect 224 276 358 288
rect 224 100 275 276
rect 332 100 358 276
rect 224 88 358 100
rect 556 88 716 288
rect 888 276 1048 288
rect 888 100 940 276
rect 996 100 1048 276
rect 888 88 1048 100
rect 1220 276 1354 289
rect 1220 100 1261 276
rect 1313 100 1354 276
rect 1220 88 1354 100
rect -36 -60 5 88
rect 1266 -60 1307 88
rect -36 -101 1307 -60
rect 260 -188 270 -136
rect 336 -188 346 -136
rect 924 -138 934 -136
rect 921 -144 934 -138
rect 921 -181 933 -144
rect 921 -187 934 -181
rect 924 -188 934 -187
rect 1000 -188 1010 -136
<< via1 >>
rect 610 889 662 941
rect 74 477 202 529
rect 74 317 202 369
rect 610 477 662 529
rect 406 317 534 369
rect 738 317 866 369
rect 1070 477 1198 529
rect 1070 317 1198 369
rect -41 100 11 276
rect 275 100 332 276
rect 940 100 996 276
rect 1261 100 1313 276
rect 270 -146 336 -136
rect 270 -180 277 -146
rect 277 -180 329 -146
rect 329 -180 336 -146
rect 270 -188 336 -180
rect 934 -144 1000 -136
rect 934 -181 998 -144
rect 998 -181 1000 -144
rect 934 -188 1000 -181
<< metal2 >>
rect 606 945 666 955
rect 606 875 666 885
rect 74 529 202 539
rect 74 448 202 477
rect 610 529 662 539
rect 1070 529 1198 539
rect 662 477 665 486
rect 610 448 665 477
rect 1070 448 1198 477
rect -41 396 1313 448
rect -41 276 11 396
rect 74 369 202 396
rect 74 307 202 317
rect 406 369 534 396
rect 406 307 534 317
rect 738 369 866 396
rect 738 307 866 317
rect 1070 369 1198 396
rect 1070 307 1198 317
rect 275 276 332 286
rect -41 90 11 100
rect 274 100 275 110
rect 274 95 332 100
rect 608 276 664 286
rect 940 276 996 286
rect 267 -60 337 95
rect 608 90 664 100
rect 934 100 940 105
rect 1261 276 1313 396
rect 996 100 1000 105
rect 934 -60 1000 100
rect 1261 90 1313 100
rect 267 -101 1000 -60
rect 267 -136 337 -101
rect 267 -167 270 -136
rect 336 -167 337 -136
rect 934 -136 1000 -101
rect 270 -198 336 -188
rect 934 -198 1000 -188
<< via2 >>
rect 606 941 666 945
rect 606 889 610 941
rect 610 889 662 941
rect 662 889 666 941
rect 606 885 666 889
rect 608 100 664 276
<< metal3 >>
rect 596 945 676 950
rect 596 885 606 945
rect 666 885 676 945
rect 596 880 676 885
rect 606 281 666 880
rect 598 276 674 281
rect 598 100 608 276
rect 664 100 674 276
rect 598 95 674 100
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_0
timestamp 1729266807
transform 1 0 -15 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_1
timestamp 1729266807
transform 1 0 -15 0 1 658
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_2
timestamp 1729266807
transform 1 0 1287 0 1 658
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_6H9P4D  sky130_fd_pr__nfet_01v8_6H9P4D_3
timestamp 1729266807
transform 1 0 1287 0 1 188
box -73 -126 73 126
use sky130_fd_pr__nfet_01v8_DB328X  sky130_fd_pr__nfet_01v8_DB328X_0
timestamp 1729266807
transform 1 0 636 0 1 658
box -636 -188 636 188
use sky130_fd_pr__nfet_01v8_DB328X  sky130_fd_pr__nfet_01v8_DB328X_1
timestamp 1729266807
transform 1 0 636 0 1 188
box -636 -188 636 188
<< labels >>
flabel metal2 963 -23 963 -23 0 FreeSans 800 0 0 0 GND
port 2 nsew
flabel metal3 635 331 635 331 0 FreeSans 800 0 0 0 OUT
port 1 nsew
flabel metal2 133 428 133 428 0 FreeSans 800 0 0 0 D6
port 0 nsew
<< end >>
