magic
tech sky130A
magscale 1 2
timestamp 1729246480
<< nwell >>
rect -176 504 622 1231
rect -176 495 281 504
rect 323 495 622 504
rect -176 -1316 622 495
<< nsubdiff >>
rect -140 1161 -80 1195
rect 526 1161 586 1195
rect -140 1135 -106 1161
rect 552 1135 586 1161
rect -140 -1246 -106 -1220
rect 552 -1246 586 -1220
rect -140 -1280 -80 -1246
rect 526 -1280 586 -1246
<< nsubdiffcont >>
rect -80 1161 526 1195
rect -140 -1220 -106 1135
rect 552 -1220 586 1135
rect -80 -1280 526 -1246
<< poly >>
rect 6 562 36 595
rect -56 546 36 562
rect -56 512 -40 546
rect -6 512 36 546
rect -56 496 36 512
rect 410 556 440 585
rect 410 540 502 556
rect 410 506 452 540
rect 486 506 502 540
rect 410 490 502 506
rect 6 68 36 90
rect -56 52 36 68
rect -56 18 -40 52
rect -6 18 36 52
rect -56 2 36 18
rect 410 69 440 96
rect 410 53 502 69
rect 410 19 452 53
rect 486 19 502 53
rect -56 -112 36 -96
rect 94 -104 194 8
rect 252 -103 352 9
rect 410 3 502 19
rect -56 -146 -40 -112
rect -6 -146 36 -112
rect -56 -162 36 -146
rect 6 -194 36 -162
rect 410 -112 502 -96
rect 410 -146 452 -112
rect 486 -146 502 -112
rect 410 -162 502 -146
rect 410 -188 440 -162
rect -56 -569 36 -553
rect -56 -603 -40 -569
rect -6 -603 36 -569
rect -56 -619 36 -603
rect 6 -680 36 -619
rect 410 -569 502 -553
rect 410 -603 452 -569
rect 486 -603 502 -569
rect 410 -619 502 -603
rect 410 -672 441 -619
<< polycont >>
rect -40 512 -6 546
rect 452 506 486 540
rect -40 18 -6 52
rect 452 19 486 53
rect -40 -146 -6 -112
rect 452 -146 486 -112
rect -40 -603 -6 -569
rect 452 -603 486 -569
<< locali >>
rect -140 1161 -80 1195
rect 526 1161 586 1195
rect -140 1135 -106 1161
rect 552 1135 586 1161
rect -40 546 -6 595
rect -56 512 -40 546
rect -6 512 10 546
rect 452 540 486 609
rect 436 506 452 540
rect 486 506 502 540
rect -40 52 -6 107
rect 452 53 486 112
rect -56 18 -40 52
rect -6 18 10 52
rect 436 19 452 53
rect 486 19 502 53
rect -56 -146 -40 -112
rect -6 -146 10 -112
rect 436 -146 452 -112
rect 486 -146 502 -112
rect -40 -200 -6 -146
rect 452 -198 486 -146
rect -56 -603 -40 -569
rect -6 -603 10 -569
rect 436 -603 452 -569
rect 486 -603 502 -569
rect -40 -693 -6 -603
rect 452 -695 486 -603
rect -140 -1246 -106 -1220
rect 552 -1246 586 -1220
rect -140 -1280 -80 -1246
rect 526 -1280 586 -1246
<< viali >>
rect 185 1161 280 1195
rect -40 512 -6 546
rect 452 506 486 540
rect -40 18 -6 52
rect 452 19 486 53
rect -40 -146 -6 -112
rect 452 -146 486 -112
rect -40 -603 -6 -569
rect 452 -603 486 -569
<< metal1 >>
rect 173 1195 292 1201
rect 173 1161 185 1195
rect 280 1161 292 1195
rect 173 1155 292 1161
rect 440 1115 446 1120
rect 0 1073 446 1115
rect 0 794 42 1073
rect 440 1068 446 1073
rect 498 1068 504 1120
rect -46 594 88 794
rect 187 606 197 782
rect 249 606 259 782
rect 358 594 399 794
rect 451 594 492 794
rect -46 552 4 594
rect -52 546 6 552
rect -52 512 -40 546
rect -6 512 6 546
rect -52 506 6 512
rect 122 465 164 513
rect 258 504 268 556
rect 336 504 346 556
rect 442 546 492 594
rect 440 540 498 546
rect 440 506 452 540
rect 486 506 498 540
rect 440 500 498 506
rect 122 423 323 465
rect 100 338 110 390
rect 178 338 188 390
rect 281 371 323 423
rect -46 288 88 300
rect 358 288 492 300
rect -59 112 -49 288
rect 3 112 88 288
rect 187 112 197 288
rect 249 112 259 288
rect 358 112 443 288
rect 495 112 505 288
rect -52 100 88 112
rect 358 100 498 112
rect -52 52 6 100
rect -52 18 -40 52
rect -6 18 6 52
rect -52 12 6 18
rect 440 53 498 100
rect 440 19 452 53
rect 486 19 498 53
rect 440 13 498 19
rect -52 -112 6 -106
rect -52 -146 -40 -112
rect -6 -146 6 -112
rect -52 -194 6 -146
rect 440 -112 498 -106
rect 440 -146 452 -112
rect 486 -146 498 -112
rect 440 -194 498 -146
rect -52 -206 88 -194
rect 358 -206 498 -194
rect -59 -382 -49 -206
rect 3 -382 88 -206
rect 187 -382 197 -206
rect 249 -382 259 -206
rect 358 -382 443 -206
rect 495 -382 505 -206
rect -46 -394 88 -382
rect 358 -394 492 -382
rect 100 -484 110 -432
rect 178 -484 188 -432
rect 280 -520 321 -478
rect 123 -561 321 -520
rect -52 -569 6 -563
rect -52 -603 -40 -569
rect -6 -603 6 -569
rect -52 -688 6 -603
rect 123 -607 164 -561
rect 440 -569 498 -563
rect 258 -650 268 -598
rect 336 -650 346 -598
rect 440 -603 452 -569
rect 486 -603 498 -569
rect 440 -688 498 -603
rect -52 -698 88 -688
rect -46 -888 88 -698
rect 187 -876 197 -700
rect 249 -876 259 -700
rect 358 -888 399 -688
rect 451 -711 498 -688
rect 451 -888 492 -711
rect 4 -1148 48 -888
rect 436 -1148 442 -1144
rect 4 -1192 442 -1148
rect 436 -1196 442 -1192
rect 494 -1196 500 -1144
<< via1 >>
rect 446 1068 498 1120
rect 197 606 249 782
rect 399 594 451 794
rect 268 504 336 556
rect 110 338 178 390
rect -49 112 3 288
rect 197 112 249 288
rect 443 112 495 288
rect -49 -382 3 -206
rect 197 -382 249 -206
rect 443 -382 495 -206
rect 110 -484 178 -432
rect 268 -650 336 -598
rect 197 -876 249 -700
rect 399 -888 451 -688
rect 442 -1196 494 -1144
<< metal2 >>
rect 442 1124 502 1134
rect 442 1054 502 1064
rect -49 935 451 987
rect -49 288 3 935
rect 399 794 451 935
rect 195 782 251 792
rect 195 596 251 606
rect 399 584 451 594
rect 268 556 336 566
rect 268 479 336 504
rect 110 411 336 479
rect 110 390 178 411
rect 110 328 178 338
rect -49 -206 3 112
rect 195 288 251 298
rect 195 102 251 112
rect 441 288 497 298
rect 441 102 497 112
rect -49 -1045 3 -382
rect 195 -206 251 -196
rect 195 -392 251 -382
rect 441 -206 497 -196
rect 441 -392 497 -382
rect 110 -432 178 -422
rect 110 -507 178 -484
rect 110 -575 336 -507
rect 268 -598 336 -575
rect 268 -660 336 -650
rect 399 -688 451 -678
rect 195 -700 251 -690
rect 195 -886 251 -876
rect 399 -1045 451 -888
rect -49 -1097 451 -1045
rect 433 -1135 503 -1125
rect 433 -1215 503 -1205
<< via2 >>
rect 442 1120 502 1124
rect 442 1068 446 1120
rect 446 1068 498 1120
rect 498 1068 502 1120
rect 442 1064 502 1068
rect 195 606 197 782
rect 197 606 249 782
rect 249 606 251 782
rect 195 112 197 288
rect 197 112 249 288
rect 249 112 251 288
rect 441 112 443 288
rect 443 112 495 288
rect 495 112 497 288
rect 195 -382 197 -206
rect 197 -382 249 -206
rect 249 -382 251 -206
rect 441 -382 443 -206
rect 443 -382 495 -206
rect 495 -382 497 -206
rect 195 -876 197 -700
rect 197 -876 249 -700
rect 249 -876 251 -700
rect 433 -1144 503 -1135
rect 433 -1196 442 -1144
rect 442 -1196 494 -1144
rect 494 -1196 503 -1144
rect 433 -1205 503 -1196
<< metal3 >>
rect 432 1124 512 1129
rect 432 1064 442 1124
rect 502 1064 512 1124
rect 432 1059 512 1064
rect 185 782 261 787
rect 185 606 195 782
rect 251 606 261 782
rect 185 601 261 606
rect 194 293 254 601
rect 442 293 504 1059
rect 185 288 261 293
rect 185 112 195 288
rect 251 112 261 288
rect 185 107 261 112
rect 431 288 507 293
rect 431 112 441 288
rect 497 112 507 288
rect 431 107 507 112
rect 194 -201 254 107
rect 442 -201 504 107
rect 185 -206 261 -201
rect 185 -382 195 -206
rect 251 -382 261 -206
rect 185 -387 261 -382
rect 431 -206 507 -201
rect 431 -382 441 -206
rect 497 -382 507 -206
rect 431 -387 507 -382
rect 194 -695 254 -387
rect 185 -700 261 -695
rect 185 -876 195 -700
rect 251 -876 261 -700
rect 185 -881 261 -876
rect 442 -1130 504 -387
rect 423 -1135 513 -1130
rect 423 -1205 433 -1135
rect 503 -1205 513 -1135
rect 423 -1210 513 -1205
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_0
timestamp 1729235383
transform 1 0 425 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_1
timestamp 1729235383
transform 1 0 21 0 1 200
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_2
timestamp 1729235383
transform 1 0 425 0 1 -788
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_3
timestamp 1729235383
transform 1 0 21 0 1 -788
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_4
timestamp 1729235383
transform 1 0 21 0 1 -294
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_5
timestamp 1729235383
transform 1 0 425 0 1 -294
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_6
timestamp 1729235383
transform 1 0 21 0 1 694
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_2XUZHN  sky130_fd_pr__pfet_01v8_2XUZHN_7
timestamp 1729235383
transform 1 0 425 0 1 694
box -109 -162 109 162
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_0
timestamp 1729235383
transform 1 0 223 0 1 -788
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_1
timestamp 1729235383
transform 1 0 223 0 1 200
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_2
timestamp 1729235383
transform 1 0 223 0 1 694
box -223 -200 223 200
use sky130_fd_pr__pfet_01v8_BHVYY6  sky130_fd_pr__pfet_01v8_BHVYY6_3
timestamp 1729235383
transform 1 0 223 0 1 -294
box -223 -200 223 200
<< labels >>
flabel viali 222 1177 222 1177 0 FreeSans 800 0 0 0 VDD
port 0 nsew
flabel metal2 123 959 123 959 0 FreeSans 800 0 0 0 D6
port 1 nsew
flabel metal3 469 1013 469 1013 0 FreeSans 800 0 0 0 OUT
port 2 nsew
flabel metal1 142 491 142 491 0 FreeSans 800 0 0 0 VIP
port 3 nsew
flabel metal3 221 318 221 318 0 FreeSans 800 0 0 0 D5
port 4 nsew
flabel metal2 301 -577 301 -577 0 FreeSans 800 0 0 0 VIN
port 5 nsew
<< end >>
