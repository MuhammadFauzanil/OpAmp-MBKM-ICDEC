magic
tech sky130A
timestamp 1729266807
<< nmos >>
rect -289 -50 -209 50
rect -123 -50 -43 50
rect 43 -50 123 50
rect 209 -50 289 50
<< ndiff >>
rect -318 44 -289 50
rect -318 -44 -312 44
rect -295 -44 -289 44
rect -318 -50 -289 -44
rect -209 44 -180 50
rect -209 -44 -203 44
rect -186 -44 -180 44
rect -209 -50 -180 -44
rect -152 44 -123 50
rect -152 -44 -146 44
rect -129 -44 -123 44
rect -152 -50 -123 -44
rect -43 44 -14 50
rect -43 -44 -37 44
rect -20 -44 -14 44
rect -43 -50 -14 -44
rect 14 44 43 50
rect 14 -44 20 44
rect 37 -44 43 44
rect 14 -50 43 -44
rect 123 44 152 50
rect 123 -44 129 44
rect 146 -44 152 44
rect 123 -50 152 -44
rect 180 44 209 50
rect 180 -44 186 44
rect 203 -44 209 44
rect 180 -50 209 -44
rect 289 44 318 50
rect 289 -44 295 44
rect 312 -44 318 44
rect 289 -50 318 -44
<< ndiffc >>
rect -312 -44 -295 44
rect -203 -44 -186 44
rect -146 -44 -129 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 129 -44 146 44
rect 186 -44 203 44
rect 295 -44 312 44
<< poly >>
rect -289 86 -209 94
rect -289 69 -281 86
rect -217 69 -209 86
rect -289 50 -209 69
rect -123 86 -43 94
rect -123 69 -115 86
rect -51 69 -43 86
rect -123 50 -43 69
rect 43 86 123 94
rect 43 69 51 86
rect 115 69 123 86
rect 43 50 123 69
rect 209 86 289 94
rect 209 69 217 86
rect 281 69 289 86
rect 209 50 289 69
rect -289 -69 -209 -50
rect -289 -86 -281 -69
rect -217 -86 -209 -69
rect -289 -94 -209 -86
rect -123 -69 -43 -50
rect -123 -86 -115 -69
rect -51 -86 -43 -69
rect -123 -94 -43 -86
rect 43 -69 123 -50
rect 43 -86 51 -69
rect 115 -86 123 -69
rect 43 -94 123 -86
rect 209 -69 289 -50
rect 209 -86 217 -69
rect 281 -86 289 -69
rect 209 -94 289 -86
<< polycont >>
rect -281 69 -217 86
rect -115 69 -51 86
rect 51 69 115 86
rect 217 69 281 86
rect -281 -86 -217 -69
rect -115 -86 -51 -69
rect 51 -86 115 -69
rect 217 -86 281 -69
<< locali >>
rect -289 69 -281 86
rect -217 69 -209 86
rect -123 69 -115 86
rect -51 69 -43 86
rect 43 69 51 86
rect 115 69 123 86
rect 209 69 217 86
rect 281 69 289 86
rect -312 44 -295 52
rect -312 -52 -295 -44
rect -203 44 -186 52
rect -203 -52 -186 -44
rect -146 44 -129 52
rect -146 -52 -129 -44
rect -37 44 -20 52
rect -37 -52 -20 -44
rect 20 44 37 52
rect 20 -52 37 -44
rect 129 44 146 52
rect 129 -52 146 -44
rect 186 44 203 52
rect 186 -52 203 -44
rect 295 44 312 52
rect 295 -52 312 -44
rect -289 -86 -281 -69
rect -217 -86 -209 -69
rect -123 -86 -115 -69
rect -51 -86 -43 -69
rect 43 -86 51 -69
rect 115 -86 123 -69
rect 209 -86 217 -69
rect 281 -86 289 -69
<< viali >>
rect -281 69 -217 86
rect -115 69 -51 86
rect 51 69 115 86
rect 217 69 281 86
rect -312 -44 -295 44
rect -203 -44 -186 44
rect -146 -44 -129 44
rect -37 -44 -20 44
rect 20 -44 37 44
rect 129 -44 146 44
rect 186 -44 203 44
rect 295 -44 312 44
rect -281 -86 -217 -69
rect -115 -86 -51 -69
rect 51 -86 115 -69
rect 217 -86 281 -69
<< metal1 >>
rect -287 86 -211 89
rect -287 69 -281 86
rect -217 69 -211 86
rect -287 66 -211 69
rect -121 86 -45 89
rect -121 69 -115 86
rect -51 69 -45 86
rect -121 66 -45 69
rect 45 86 121 89
rect 45 69 51 86
rect 115 69 121 86
rect 45 66 121 69
rect 211 86 287 89
rect 211 69 217 86
rect 281 69 287 86
rect 211 66 287 69
rect -315 44 -292 50
rect -315 -44 -312 44
rect -295 -44 -292 44
rect -315 -50 -292 -44
rect -206 44 -183 50
rect -206 -44 -203 44
rect -186 -44 -183 44
rect -206 -50 -183 -44
rect -149 44 -126 50
rect -149 -44 -146 44
rect -129 -44 -126 44
rect -149 -50 -126 -44
rect -40 44 -17 50
rect -40 -44 -37 44
rect -20 -44 -17 44
rect -40 -50 -17 -44
rect 17 44 40 50
rect 17 -44 20 44
rect 37 -44 40 44
rect 17 -50 40 -44
rect 126 44 149 50
rect 126 -44 129 44
rect 146 -44 149 44
rect 126 -50 149 -44
rect 183 44 206 50
rect 183 -44 186 44
rect 203 -44 206 44
rect 183 -50 206 -44
rect 292 44 315 50
rect 292 -44 295 44
rect 312 -44 315 44
rect 292 -50 315 -44
rect -287 -69 -211 -66
rect -287 -86 -281 -69
rect -217 -86 -211 -69
rect -287 -89 -211 -86
rect -121 -69 -45 -66
rect -121 -86 -115 -69
rect -51 -86 -45 -69
rect -121 -89 -45 -86
rect 45 -69 121 -66
rect 45 -86 51 -69
rect 115 -86 121 -69
rect 45 -89 121 -86
rect 211 -69 287 -66
rect 211 -86 217 -69
rect 281 -86 287 -69
rect 211 -89 287 -86
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 1 nf 4 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
